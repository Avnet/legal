------------------------------------------------------------------------------
--      _____
--     *     *
--    *____   *____
--   * *===*   *==*
--  *___*===*___**  AVNET
--       *======*
--        *====*
------------------------------------------------------------------------------
--
-- This design is the property of Avnet.  Publication of this
-- design is not authorized without written consent from Avnet.
--
-- Please direct any questions to the Avnet Technical Community:
--    http://community.em.avnet.com/
--
-- Product information is available at:
--    http://www.em.avnet.com/arty
--
-- Disclaimer:
--    Avnet, Inc. makes no warranty for the use of this code or design.
--    This code is provided  "As Is". Avnet, Inc assumes no responsibility for
--    any errors, which may appear in this code, nor does it make a commitment
--    to update the information contained herein. Avnet, Inc specifically
--    disclaims any implied warranties of fitness for a particular purpose.
--                     Copyright(c) 2015 Avnet, Inc.
--                             All rights reserved.
--
------------------------------------------------------------------------------
--
-- Create Date:         Aug 09, 2015
-- Design Name:         MAX44000 Example Application
-- Module Name:         MAX44000.vhd
-- Project Name:        Arty Example Code
-- Target Devices:      Xilinx Artix-7 35T
-- Hardware Boards:     Arty, Maxim MAX44000PMB1 Pmod
--
-- Tool versions:       Xilinx Vivado 2015.2
--
-- Description:         This example reads the ambient light using the 
--                      Maxim MAX44000PMB1 Pmod
--
-- Dependencies:
--
-- Revision:            Aug 09, 2015: 1.00 Initial version
--
------------------------------------------------------------------------------
