------------------------------------------------------------------------------
--      _____
--     *     *
--    *____   *____
--   * *===*   *==*
--  *___*===*___**  AVNET
--       *======*
--        *====*
------------------------------------------------------------------------------
--
-- This design is the property of Avnet.  Publication of this
-- design is not authorized without written consent from Avnet.
--
-- Please direct any questions to the PicoZed community support forum:
--    http://www.picozed.org/forum
--
-- Product information is available at:
--    http://www.picozed.org/product/picozed
--
-- Disclaimer:
--    Avnet, Inc. makes no warranty for the use of this code or design.
--    This code is provided  "As Is". Avnet, Inc assumes no responsibility for
--    any errors, which may appear in this code, nor does it make a commitment
--    to update the information contained herein. Avnet, Inc specifically
--    disclaims any implied warranties of fitness for a particular purpose.
--                     Copyright(c) 2016 Avnet, Inc.
--                             All rights reserved.
--
------------------------------------------------------------------------------
--
-- Create Date:         Nov 10, 2015
-- Design Name:         PicoZed FMC2 Carrier MAC ID Test
-- Module Name:         unio_eeprom_test.vhd
-- Project Name:        PicoZed FMC2 Carrier MAC ID Test
-- Target Devices:      Xilinx Zynq-7000
-- Hardware Boards:     PicoZed, PicoZed FMC2 Carrier
--
-- Tool versions:       Xilinx Vivado 2015.2
--
-- Description:         Microchip UNI/O EEPROM test for PicoZed FMC2 Carrier
--
-- Dependencies:
--
-- Revision:            Nov 10, 2015: 1.00 Initial version
--
------------------------------------------------------------------------------
